// map_colorizer.v
// Thong & Deepen
//
// Determine color at a given map position, based on the pixel position and map value

module map_colorizer
#(
  parameter COLOR_WIDTH = 12,
  parameter SPRITE_BLACK = 0,
  parameter SPRITE_WALL  = 0,
  parameter SPRITE_EMPTY = 0
)(
  input wire [1:0]       map_value,      // map value returned from the map memory
  input wire [11:0]      pixel_row,      // pixel row from the dtg
  input wire [11:0]      pixel_column,   // pixel column from the dtg
  input wire             out_of_map,     // indicate if the given pixel coordinates is out of the map (1) or not (0)
  output reg [11:0] map_color  
);

// ==================================================
// DECLARATIONS
// ==================================================

// adjust map value based on the out_of_map signal
wire [1:0] map_value_adjusted;

// sand sprite
reg [767:0] sprite_sand = {
  12'h7b9,
  12'hca6,
  12'hc95,
  12'hc95,
  12'hc95,
  12'hca6,
  12'hc95,
  12'h7b9,
  12'hed9,
  12'hdc8,
  12'hed9,
  12'hdc8,
  12'hca6,
  12'hdc8,
  12'hdc8,
  12'hc95,
  12'hc95,
  12'hca6,
  12'hdc8,
  12'hca6,
  12'hdc8,
  12'hca6,
  12'hdc8,
  12'hed9,
  12'hca6,
  12'hdc8,
  12'hdc8,
  12'hdc8,
  12'hed9,
  12'hdc8,
  12'hdc8,
  12'hca6,
  12'hc95,
  12'hca6,
  12'hdc8,
  12'hca6,
  12'hdc8,
  12'hdc8,
  12'hdc8,
  12'hc95,
  12'hca6,
  12'hdc8,
  12'hdc8,
  12'hdc8,
  12'hdc8,
  12'hdc8,
  12'hca6,
  12'hc95,
  12'hc95,
  12'hdc8,
  12'hdc8,
  12'hdc8,
  12'hdc8,
  12'hdc8,
  12'hdc8,
  12'hc95,
  12'h7b9,
  12'hc95,
  12'hc95,
  12'hed9,
  12'hc95,
  12'hca6,
  12'hc95,
  12'h7b9
};

// grass sprite - changed to solid sky color
reg [767:0] sprite_grass = {
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e,
  12'h58e
};

// road sprite - changed to bandicoot road
reg [3071:0] sprite_road = {
  12'h8b0,
  12'h8b0,
  12'h8b0,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h8b0,
  12'h8b0,
  12'h8b0,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h680,
  12'h680,
  12'h8b0,
  12'h680,
  12'h680,
  12'h690,
  12'h690,
  12'h680,
  12'h680,
  12'h690,
  12'h8b0,
  12'h690,
  12'h680,
  12'h680,
  12'h690,
  12'h690,
  12'h680,
  12'h680,
  12'h570,
  12'h570,
  12'h570,
  12'h680,
  12'h680,
  12'h570,
  12'h570,
  12'h680,
  12'h690,
  12'h680,
  12'h570,
  12'h570,
  12'h570,
  12'h570,
  12'h680,
  12'hb81,
  12'hb81,
  12'hb81,
  12'hb81,
  12'hb81,
  12'h570,
  12'h570,
  12'hb81,
  12'h570,
  12'h570,
  12'h570,
  12'h570,
  12'hb81,
  12'hb81,
  12'hb81,
  12'h570,
  12'hc90,
  12'hda0,
  12'hc90,
  12'hc90,
  12'hc90,
  12'hda0,
  12'hda0,
  12'hda0,
  12'h570,
  12'h570,
  12'hc90,
  12'hc90,
  12'hda0,
  12'hda0,
  12'hc90,
  12'hc90,
  12'heb0,
  12'heb0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hda0,
  12'hda0,
  12'heb0,
  12'heb0,
  12'heb0,
  12'heb0,
  12'heb0,
  12'heb0,
  12'heb0,
  12'heb0,
  12'heb0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfe8,
  12'hfe8,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hda0,
  12'hda0,
  12'heb0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfd4,
  12'hfd4,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'heb0,
  12'hfc0,
  12'hfd4,
  12'hfe8,
  12'hfe8,
  12'hfd4,
  12'hfc0,
  12'hfc0,
  12'heb0,
  12'heb0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'hfc0,
  12'heb0,
  12'heb0,
  12'h680,
  12'hda0,
  12'hda0,
  12'hda0,
  12'h690,
  12'hda0,
  12'hda0,
  12'hda0,
  12'hda0,
  12'hda0,
  12'hda0,
  12'hda0,
  12'hda0,
  12'hda0,
  12'hda0,
  12'h690,
  12'h8b0,
  12'h680,
  12'hda0,
  12'h690,
  12'h8b0,
  12'h690,
  12'hda0,
  12'h680,
  12'h690,
  12'h690,
  12'hda0,
  12'h690,
  12'h690,
  12'hda0,
  12'h690,
  12'h8b0,
  12'h8b0,
  12'h8b0,
  12'h690,
  12'h8b0,
  12'h8b0,
  12'h8b0,
  12'h680,
  12'h680,
  12'h8b0,
  12'h8b0,
  12'h690,
  12'h690,
  12'h8b0,
  12'h690,
  12'h690,
  12'h8b0,
  12'h690,
  12'h690,
  12'h690,
  12'h8b0,
  12'h8b0,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h690,
  12'h680,
  12'h680,
  12'h450,
  12'h450,
  12'h570,
  12'h570,
  12'h690,
  12'h690,
  12'h570,
  12'h690,
  12'h690,
  12'h680,
  12'h570,
  12'h680,
  12'h570,
  12'h450,
  12'h450,
  12'h450,
  12'h521,
  12'h521,
  12'h521,
  12'h570,
  12'h570,
  12'h450,
  12'h570,
  12'h570,
  12'h570,
  12'h450,
  12'h450,
  12'h521,
  12'h521,
  12'h521,
  12'h521,
  12'h521,
  12'h521,
  12'h521,
  12'h521,
  12'h521,
  12'h450,
  12'h450,
  12'h521,
  12'h450,
  12'h450,
  12'h521,
  12'h521
};

// flower sprite
reg [767:0] sprite_flower = {
  12'h420,
  12'h420,
  12'h520,
  12'h520,
  12'h520,
  12'h520,
  12'h631,
  12'h631,
  12'h420,
  12'h620,
  12'h620,
  12'h420,
  12'h520,
  12'h520,
  12'h520,
  12'h631,
  12'h420,
  12'h630,
  12'h420,
  12'h520,
  12'h420,
  12'h520,
  12'h520,
  12'h520,
  12'h420,
  12'h420,
  12'h520,
  12'h520,
  12'h520,
  12'h420,
  12'h420,
  12'h731,
  12'h420,
  12'h520,
  12'h520,
  12'h520,
  12'h520,
  12'h520,
  12'h420,
  12'h741,
  12'h420,
  12'h420,
  12'h620,
  12'h520,
  12'h520,
  12'h520,
  12'h520,
  12'h530,
  12'h420,
  12'h420,
  12'h420,
  12'h620,
  12'h520,
  12'h520,
  12'h420,
  12'h520,
  12'h420,
  12'h630,
  12'h420,
  12'h420,
  12'h420,
  12'h520,
  12'h520,
  12'h520
};

// ==================================================
// LOGIC
// ==================================================

// adjust map value to '00 (empty) if current pixel is out of the map
assign map_value_adjusted = out_of_map ? 2'b00 : map_value;

// determine color based on map value
always @(*) begin
  map_color = 12'h000;
  case (map_value_adjusted)
    2'b00: map_color = sprite_grass [(12'd63 -  ((pixel_row[2:0] << 3) +  pixel_column[2:0]))*12+:12 ];
    2'b01: map_color = sprite_road  [(12'd255 - ((pixel_row[3:0] << 4) +  pixel_column[3:0]))*12+:12 ];
    2'b10: map_color = sprite_flower[(12'd63 -  ((pixel_row[2:0] << 3) +  pixel_column[2:0]))*12+:12 ];
    default: map_color = 12'h000;
  endcase
end

endmodule